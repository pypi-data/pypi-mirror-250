*
.SUBCKT newckt a b c
* new subckt
R a b 1k
C b c 1pF
.ENDS
